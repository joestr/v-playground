module main

/*
	Using the println() function to print a text on the screen
*/
fn main() {
	println('testing out vlang') // try replacing the single quotes (') with double quotes (")
}