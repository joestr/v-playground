module main

/*
	Intialize two integer variables and print out.

	Add them both together and print them out in the form of 'Result: x' (replace x with the result)
*/
fn main() {
	a := 1 // assign variables with :=
	b := 2
	println(a)
	println(b)
	c := a + b
	println("Result: $c")
}