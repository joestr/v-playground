module main

fn main() {
	println('testing out vlang')
}